.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}

vds common gnd 0
vgs gate gnd 1.8
vdum1 common drain1 0
vdum2 common drain2 0 

M1      drain1       gate     drain2     drain2  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2     drain2       gate       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M3      drain1       gate       gnd     gnd  CMOSN   W={width_N}   L={2*2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.dc vds 0 1.8 0.01 

.control 
run 
plot (vdum1#branch) (vdum2#branch) vs v(common)
.endc